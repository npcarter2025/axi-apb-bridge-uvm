`ifndef APB_SEQUENCER_SVH
`define APB_SEQUENCER_SVH

typedef uvm_sequencer #(apb_transaction) apb_sequencer;

`endif

