

interface axi_lite_if;


endinterface