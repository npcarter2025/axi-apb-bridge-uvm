`ifndef AXI_LITE_SEQUENCER_SVH
`define AXI_LITE_SEQUENCER_SVH

typedef uvm_sequencer #(axi_lite_transaction) axi_lite_sequencer;

`endif
